module Train_Display_Generator(clock,act_D,addr16[15:0],disp10[9:0]);
	
	// PI and PO
	input act_D;
	input clock;
	input [15:0] addr16;	
	
	output [9:0] disp10; 
	
	reg [9:0] disp10;
	
always @(posedge clock)
	if(act_D == 1) begin
		case(addr16)

		16'b0000000000000000: disp10 <= 10'b0000000000;
		16'b0000000100100011: disp10 <= 10'b0000001111;
		16'b0001001000110100: disp10 <= 10'b0000011110;
		16'b0010001101000101: disp10 <= 10'b0000111100;
		16'b0011010001010110: disp10 <= 10'b0001111000;
		16'b0100010101100111: disp10 <= 10'b0011110000;
		16'b0101011001111000: disp10 <= 10'b0111100000;
		16'b0110011110001001: disp10 <= 10'b1111000000;
		//16'b01111000: disp10 <= 10'b0110000000;
		//16'b10001001: disp10 <= 10'b1100000000;
		16'b0000000011111111: disp10 <= 10'b0000000000;
		16'b0000000111111111: disp10 <= 10'b0000000011;
		16'b0001001011111111: disp10 <= 10'b0000000110;
		16'b0010001111111111: disp10 <= 10'b0000001100;
		16'b0011010011111111: disp10 <= 10'b0000011000;
		16'b0100010111111111: disp10 <= 10'b0000110000;
		16'b0101011011111111: disp10 <= 10'b0001100000;
		16'b0110011111111111: disp10 <= 10'b0011000000;
		16'b0111100011111111: disp10 <= 10'b0110000000;
		16'b1000100111111111: disp10 <= 10'b1100000000;		
		
		default:	disp10 <= 10'b0000000000;  // Number other than 0-9 is not displayed 

		endcase
	end
	else begin
		disp10 <= 10'b0000000000;
	end	
endmodule
